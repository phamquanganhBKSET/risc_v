`define INST_WIDTH      32
`define REG_WIDTH       32
`define NUM_REG         32
`define MEM_WIDTH       8
`define IMM_WIDTH       12
`define IMM_WIDTH_U     20
`define IMEM_DEPTH      2**10 // 1KB
`define DMEM_DEPTH      2**20 // 1MB
`define REG_ADDR_WIDTH  $clog2(NUM_REG)
`define PC_WIDTH        $clog2(IMEM_DEPTH)
`define DMEM_ADDR_WIDTH $clog2(DMEM_DEPTH)
`define IMM_SEL_I       2'b00
`define IMM_SEL_S       2'b01
`define IMM_SEL_B       2'b10
`define IMM_SEL_U       2'b11
`define IMM_SEL_WIDTH   2
`define ADD             5'b0110011
`define ADD_FUNCT3      3'h0
`define ADD_FUNCT7      7'h00
`define SUB             5'b0110011
`define SUB_FUNCT3      3'h0
`define SUB_FUNCT7      7'h20
`define XOR             5'b0110011
`define XOR_FUNCT3      3'h4
`define XOR_FUNCT7      7'h00
`define OR              5'b0110011
`define OR_FUNCT3       3'h6
`define OR_FUNCT7       7'h00
`define AND             5'b0110011
`define AND_FUNCT3      3'h7
`define AND_FUNCT7      7'h00
`define SLL             5'b0110011
`define SLL_FUNCT3      3'h1
`define SLL_FUNCT7      7'h00
`define SRL             5'b0110011
`define SRL_FUNCT3      3'h5
`define SRL_FUNCT7      7'h00
`define SRA             5'b0110011
`define SRA_FUNCT3      3'h5
`define SRA_FUNCT7      7'h20
`define SLT             5'b0110011
`define SLT_FUNCT3      3'h2
`define SLT_FUNCT7      7'h00
`define SLTU            5'b0110011
`define SLTU_FUNCT3     3'h3
`define SLTU_FUNCT7     7'h00
`define ADDI            5'b0010011
`define ADDI_FUNCT3     3'h0
`define XORI            5'b0010011
`define XORI_FUNCT3     3'h4
`define ORI             5'b0010011
`define ORI_FUNCT3      3'h6
`define ANDI            5'b0010011
`define ANDI_FUNCT3     3'h7
`define SLLI            5'b0010011
`define SLLI_FUNCT3     3'h1
`define SLLI_FUNCT7     7'h00
`define SRLI            5'b0010011
`define SRLI_FUNCT3     3'h5
`define SRLI_FUNCT7     7'h00
`define SRAI            5'b0010011
`define SRAI_FUNCT3     3'h5
`define SRAI_FUNCT7     7'h20
`define SLTI            5'b0010011
`define SLTI_FUNCT3     3'h2
`define SLTIU           5'b0010011
`define SLTIU_FUNCT3    3'h3
`define LB              5'b0000011
`define LB_FUNCT3       3'h0
`define LH              5'b0000011
`define LH_FUNCT3       3'h1
`define LW              5'b0000011
`define LW_FUNCT3       3'h2
`define LBU             5'b0000011
`define LBU_FUNCT3      3'h4
`define LHU             5'b0000011
`define LHU_FUNCT3      3'h5
`define SB              5'b0100011
`define SB_FUNCT3       3'h0
`define SH              5'b0100011
`define SH_FUNCT3       3'h1
`define SW              5'b0100011
`define SW_FUNCT3       3'h2
`define BEQ             5'b1100111
`define BEQ_FUNCT3      3'h0
`define BNE             5'b1100111
`define BNE_FUNCT3      3'h1
`define BLT             5'b1100111
`define BLT_FUNCT3      3'h4
`define BGE             5'b1100111
`define BGE_FUNCT3      3'h5
`define BLTU            5'b1100111
`define BLTU_FUNCT3     3'h6
`define BGEU            5'b1100111
`define BGEU_FUNCT3     3'h7
`define JAL             5'b1101111
`define JALR            5'b1100111
`define JALR_FUNCT3     3'h0
`define LUI             5'b0110111
`define AUIPC           5'b0010111
`define ECALL           5'b1110011
`define ECALL_FUNCT3    3'h0
`define EBREAK          5'b1110011
`define EBREAK_FUNCT3   3'h0
