`define INST_WIDTH      32
`define REG_WIDTH       5'd32
`define NUM_REG         32
`define MEM_WIDTH       8
`define IMM_WIDTH       12
`define IMM_WIDTH_U     20
`define IMEM_DEPTH      2**10 // 1KB
`define DMEM_DEPTH      2**20 // 1MB
`define REG_ADDR_WIDTH  $clog2(`NUM_REG)
`define PC_WIDTH        $clog2(`IMEM_DEPTH)
`define DMEM_ADDR_WIDTH $clog2(`DMEM_DEPTH)
`define IMM_SEL_I       2'b00
`define IMM_SEL_S       2'b01
`define IMM_SEL_B       2'b10
`define IMM_SEL_J       2'b11
`define IMM_SEL_WIDTH   2
`define ADD             7'b0110011
`define ADD_FUNCT3      3'h0
`define ADD_FUNCT7      7'h00
`define SUB             7'b0110011
`define SUB_FUNCT3      3'h0
`define SUB_FUNCT7      7'h20
`define XOR             7'b0110011
`define XOR_FUNCT3      3'h4
`define XOR_FUNCT7      7'h00
`define OR              7'b0110011
`define OR_FUNCT3       3'h6
`define OR_FUNCT7       7'h00
`define AND             7'b0110011
`define AND_FUNCT3      3'h7
`define AND_FUNCT7      7'h00
`define SLL             7'b0110011
`define SLL_FUNCT3      3'h1
`define SLL_FUNCT7      7'h00
`define SRL             7'b0110011
`define SRL_FUNCT3      3'h5
`define SRL_FUNCT7      7'h00
`define SRA             7'b0110011
`define SRA_FUNCT3      3'h5
`define SRA_FUNCT7      7'h20
`define SLT             7'b0110011
`define SLT_FUNCT3      3'h2
`define SLT_FUNCT7      7'h00
`define SLTU            7'b0110011
`define SLTU_FUNCT3     3'h3
`define SLTU_FUNCT7     7'h00
`define ADDI            7'b0010011
`define ADDI_FUNCT3     3'h0
`define XORI            7'b0010011
`define XORI_FUNCT3     3'h4
`define ORI             7'b0010011
`define ORI_FUNCT3      3'h6
`define ANDI            7'b0010011
`define ANDI_FUNCT3     3'h7
`define SLLI            7'b0010011
`define SLLI_FUNCT3     3'h1
`define SLLI_FUNCT7     7'h00
`define SRLI            7'b0010011
`define SRLI_FUNCT3     3'h5
`define SRLI_FUNCT7     7'h00
`define SRAI            7'b0010011
`define SRAI_FUNCT3     3'h5
`define SRAI_FUNCT7     7'h20
`define SLTI            7'b0010011
`define SLTI_FUNCT3     3'h2
`define SLTIU           7'b0010011
`define SLTIU_FUNCT3    3'h3
`define LB              7'b0000011
`define LB_FUNCT3       3'h0
`define LH              7'b0000011
`define LH_FUNCT3       3'h1
`define LW              7'b0000011
`define LW_FUNCT3       3'h2
`define LBU             7'b0000011
`define LBU_FUNCT3      3'h4
`define LHU             7'b0000011
`define LHU_FUNCT3      3'h5
`define SB              7'b0100011
`define SB_FUNCT3       3'h0
`define SH              7'b0100011
`define SH_FUNCT3       3'h1
`define SW              7'b0100011
`define SW_FUNCT3       3'h2
`define BEQ             7'b1100111
`define BEQ_FUNCT3      3'h0
`define BNE             7'b1100111
`define BNE_FUNCT3      3'h1
`define BLT             7'b1100111
`define BLT_FUNCT3      3'h4
`define BGE             7'b1100111
`define BGE_FUNCT3      3'h5
`define BLTU            7'b1100111
`define BLTU_FUNCT3     3'h6
`define BGEU            7'b1100111
`define BGEU_FUNCT3     3'h7
`define JAL             7'b1101111
`define JALR            7'b1100111
`define JALR_FUNCT3     3'h0
`define LUI             7'b0110111
`define AUIPC           7'b0010111
`define ECALL           7'b1110011
`define ECALL_FUNCT3    3'h0
`define EBREAK          7'b1110011
`define EBREAK_FUNCT3   3'h0
